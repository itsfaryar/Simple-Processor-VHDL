entity Memory is
end Memory;

--}} End of automatically maintained section

architecture Memory of Memory is
begin

	 -- enter your statements here --

end Memory;
